module decoder(
    input _CR,
    input [31:0] display_time,
    input [7:0] index,
    input adjust,
    input CP_1KHz,
    output [7:0] select_light,
    output [7:0] display_char
    );
endmodule
