module counter_sec(
    input CP_1Hz,
    input adjust,
    input _CR,
    input mode,
    input PE,
    input [7:0] pre_sec,
    output [7:0] show_sec,
    output cin_sec
    );
endmodule
