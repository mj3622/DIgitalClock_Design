module counter_hour(
    input cin_min,
    input PE,
    input _CR,
    input [7:0] pre_hour,
    output [7:0] show_hour,
    output cin_hour
    );
endmodule
