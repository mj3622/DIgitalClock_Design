module counter_min(
    input cin_sec,
    input [7:0] pre_min,
    input _CR,
    input PE,
    output cin_min,
    output [7:0] show_min
    );
endmodule
