module reminder(
    input _CR,
    input CP_1Hz,
    input start_light_hour,
    input start_light_alarm,
    input show_hour,
    output [15:0] start_light
);

endmodule