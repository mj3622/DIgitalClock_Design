module splitter(
    input _CR,
    input [31:0] display_time,
    input time_mode,
    input mode,
    output [7:0] pre_sec,
    output [7:0] pre_min,
    output [7:0] pre_hour,
    output PE_alarm,
    output PE_counter
    );
endmodule
